package shared_pkg;

	bit test_finished;
	int correct_count = 0, error_count = 0;
	
endpackage : shared_pkg